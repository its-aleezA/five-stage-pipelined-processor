module ControlUnit(
    input [5:0] opcode,
	 input [5:0] func,
	 output reg memtoreg,
	 output reg memwrite,
	 output reg branch,
	 output reg [2:0] aluControl,
	 output reg aluSrc,
	 output reg regdst,
	 output reg regwrite,
	 output reg jump,
	 output reg memRead
    );
	 
	 always@(opcode or func)
	 begin
	 case(opcode)
	 ///xori
	 6'b001001:
	 begin
	 aluControl<=3'b111;
	 memtoreg<=0;
	 branch<=1'b0;
	 aluSrc<=1'b1;
	 regdst<=1'b0;
	 regwrite<=1'b1;
	 jump<=1'b0;
	 memRead<=1'b0;
	 end
	 //slti
	 6'b001000:
	 begin
	 aluControl<=3'b101;
	 memtoreg<=0;
	 branch<=1'b0;
	 aluSrc<=1'b1;
	 regdst<=1'b1;
	 regwrite<=1'b1;
	 jump<=1'b0;
	 memRead<=1'b0;
	 end
	 //slt
	 6'b000111:
	 begin
	 aluControl<=3'b111;
	 memtoreg<=0;
	 branch<=1'b0;
	 aluSrc<=1'b0;
	 regdst<=1'b1;
	 regwrite<=1'b1;
	 jump<=1'b0;
	 memRead<=1'b0;
	 end
	 //and
	 6'b000110:
	 begin
	 aluControl<=3'b011;
	 memtoreg<=0;
	 branch<=1'b0;
	 aluSrc<=1'b1;
	 regdst<=1'b0;
	 regwrite<=1'b1;
	 jump<=1'b0;
	 memRead<=1'b0;
	 end
	 //lui
	 6'b000101:
	 begin
	 aluControl<=3'b010;
	 memtoreg<=2'b10;
	 branch<=1'b0;
	 aluSrc<=1'b0;
	 regdst<=1'b0;
	 regwrite<=1'b1;
	 jump<=1'b0;
	 memRead<=1'b0;
	 end
	 //lw
	 6'b000000:
	 begin
	 aluControl<=3'b010;
	 memtoreg<=1'b1;
	 branch<=1'b0;
	 aluSrc<=1'b1;
	 memwrite<=1'b0;
	 regdst<=1'b1;
	 regwrite<=1'b0;
	 jump<=1'b0;
	 memRead<=1'b1;
	 end
	 //sw
	 6'b000001:
	 begin
	 aluControl<=3'b010;
	 memtoreg<=1'b0;
	 memwrite<=1'b1;
	 branch<=1'b0;
	 aluSrc<=1'b1;
	 regdst<=1'b0;
	 regwrite<=1'b0;
	 jump<=1'b0;
	 memRead<=1'b0;
	 end
	 //beq
	 6'b000010:
	 begin
	 aluControl<=3'b110;
	 memtoreg<=1'b0;
	 memwrite<=1'b0;
	 branch<=1'b1;
	 aluSrc<=1'b0;
	 regdst<=1'b0;
	 regwrite<=1'b0;
	 jump<=1'b0;
	 memRead<=1'b0;
	 end
	 //jump
	 6'b000011:
	 begin
	 aluControl<=3'b010;
	 memtoreg<=2'b00;
	 memwrite<=1'b1;
	 branch<=1'b0;
	 aluSrc<=1'b0;
	 regdst<=1'b1;
	 regwrite<=1'b1;
	 jump<=1'b1;
	 memRead<=1'b0;
	 end
	 6'b000100:
	 case(func)
	 //add
	 6'b100000:
	 begin
	 aluControl<=3'b010;
	 memtoreg<=2'b00;
	 memwrite<=1'b1;
	 branch<=1'b0;
	 aluSrc<=1'b0;
	 regdst<=1'b1;
	 regwrite<=1'b1;
	 jump<=1'b0;
	 memRead<=1'b0;
	 end
	 //sub
	 6'b100010:
	 begin
	 aluControl<=3'b110;
	 memtoreg<=2'b00;
	 memwrite<=1'b1;
	 branch<=1'b0;
	 aluSrc<=1'b0;
	 regdst<=1'b1;
	 regwrite<=1'b1;
	 jump<=1'b0;
	 memRead<=1'b0;
	 end
	 //and
	 6'b100100:
	 begin
	 aluControl<=3'b011;
	 memtoreg<=2'b00;
	 memwrite<=1'b1;
	 branch<=1'b0;
	 aluSrc<=1'b0;
	 regdst<=1'b1;
	 regwrite<=1'b1;
	 jump<=1'b0;
	 memRead<=1'b0;
	 end
	 //or
	 6'b100101:
	 begin
	 aluControl<=3'b001;
	 memtoreg<=2'b00;
	 memwrite<=1'b1;
	 branch<=1'b0;
	 aluSrc<=1'b0;
	 regdst<=1'b1;
	 regwrite<=1'b1;
	 jump<=1'b0;
	 memRead<=1'b0;
	 end
	 //set on less than
	 6'b101010:
	 begin
	 aluControl<=3'b111;
	 memtoreg<=2'b00;
	 memwrite<=1'b1;
	 branch<=1'b0;
	 aluSrc<=1'b0;
	 regdst<=1'b1;
	 regwrite<=1'b1;
	 jump<=1'b0;
	 memRead<=1'b0;
	 end
	 default:
	 begin
	 aluControl<=3'b000;
	 memtoreg<=2'b00;
	 memwrite<=1'b0;
	 branch<=1'b0;
	 aluSrc<=1'b0;
	 regdst<=1'b0;
	 regwrite<=1'b0;
	 jump<=1'b0;
	 memRead<=1'b0;
	 end
	 endcase
	 default:
	 begin
	 aluControl<=3'b000;
	 memtoreg<=2'b00;
	 memwrite<=1'b0;
	 branch<=1'b0;
	 aluSrc<=1'b0;
	 regdst<=1'b0;
	 regwrite<=1'b0;
	 jump<=1'b0;
	 memRead<=1'b0;
	 end
	 endcase
	 end	


endmodule
