module inst_mem #(parameter N=32, D =32)(
    input [N-1:0] address,
    output reg [N-1:0] instruction
    );

	 reg [N-1:0] memory [D-1:0];
	 initial
	 begin
memory[0] = 32'b000000_00000_01001_00001_00000_000000;  // lw   $t1, 0($t0)
memory[1] = 32'b000100_00001_01011_01010_00000_100000;  // add  $t2, $t1, $t3
memory[2] = 32'b000100_01001_01011_01010_00000_100000;  // add  $t2, $t1, $t3
memory[3] = 32'b000001_00000_01001_00001_00000_000000;  // sw   $t1, 0($t0)
memory[4] = 32'b000100_01010_00001_00000_00000_100010;  // sub
memory[5] = 32'b000100_00010_00001_00000_00000_100101; // or
memory[6] = 32'b000100_00010_00001_00000_00000_100100; // and
memory[7] = 32'b000010_00101_00101_00000_00000_000001;  // beq
memory[8] = 32'b000000_00000_01001_00001_00000_000000;  // lw   $t1, 0($t0)
memory[9] = 32'b000000_00000_01001_00001_00000_000000;  // lw   $t1, 0($t0)
memory[10] = 32'b000100_00001_01011_01010_00000_100000;  // add  $t2, $t1, $t3
memory[11] = 32'b000100_01010_00001_00000_00000_100010;  // sub
memory[12] = 32'b000011_00000_00000_00000_00000_000010; // jump
memory[13] = 32'b000000_00000_01001_00001_00000_000000;  // lw   $t1, 0($t0)
memory[14] = 32'b000000_00000_01001_00001_00000_000000;  // lw   $t1, 0($t0)
memory[15] = 32'b000100_00010_00001_00000_00000_000001;
memory[16] = 32'b000001_00010_00001_00000_00000_000100;  // sw
memory[17] = 32'b000100_00010_00001_00000_00000_000001;
memory[18] = 32'b000100_00010_00001_00000_00000_000001;
memory[19] = 32'b000100_00010_00001_00000_00000_100101; // or
memory[20] = 32'b000000_00010_00001_00000_00000_000100;  // lw
memory[21] = 32'b000100_00010_00001_00000_00000_000001;
memory[22] = 32'b000100_00010_00001_00000_00000_000001;
memory[23] = 32'b000100_00010_00001_00000_00000_000001;
memory[24] = 32'b000100_00010_00001_00000_00000_000001;
memory[25] = 32'b000100_00010_00001_00000_00000_000001;
memory[26] = 32'b000100_00010_00001_00000_00000_000001;
memory[27] = 32'b000100_00010_00001_00000_00000_000001;
memory[28] = 32'b000100_00010_00001_00000_00000_000001;
memory[29] = 32'b000100_00010_00001_00000_00000_000001;
memory[30] = 32'b000100_00010_00001_00000_00000_000001;
memory[31] = 32'b000100_00010_00001_00000_00000_000001;

	 end
	 always @(address)
	 begin
	 instruction=memory[address];
	 end

endmodule
